interface ha_intf();

  logic a,b;
  logic sum,carry;
  
endinterface