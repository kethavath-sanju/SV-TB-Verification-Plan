package ha_pkg;
   
`include "ha_interface.sv"
`include "packet.sv"
`include "generator.sv"
`include "driver.sv"
`include "environment.sv"
 
 endpackage